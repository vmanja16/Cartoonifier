module tb_intensity(

);